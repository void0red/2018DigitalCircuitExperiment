-- hps.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity hps is
	port (
		clk_clk            : in    std_logic                     := '0';             --    clk.clk
		memory_mem_a       : out   std_logic_vector(12 downto 0);                    -- memory.mem_a
		memory_mem_ba      : out   std_logic_vector(2 downto 0);                     --       .mem_ba
		memory_mem_ck      : out   std_logic;                                        --       .mem_ck
		memory_mem_ck_n    : out   std_logic;                                        --       .mem_ck_n
		memory_mem_cke     : out   std_logic;                                        --       .mem_cke
		memory_mem_cs_n    : out   std_logic;                                        --       .mem_cs_n
		memory_mem_ras_n   : out   std_logic;                                        --       .mem_ras_n
		memory_mem_cas_n   : out   std_logic;                                        --       .mem_cas_n
		memory_mem_we_n    : out   std_logic;                                        --       .mem_we_n
		memory_mem_reset_n : out   std_logic;                                        --       .mem_reset_n
		memory_mem_dq      : inout std_logic_vector(7 downto 0)  := (others => '0'); --       .mem_dq
		memory_mem_dqs     : inout std_logic                     := '0';             --       .mem_dqs
		memory_mem_dqs_n   : inout std_logic                     := '0';             --       .mem_dqs_n
		memory_mem_odt     : out   std_logic;                                        --       .mem_odt
		memory_mem_dm      : out   std_logic;                                        --       .mem_dm
		memory_oct_rzqin   : in    std_logic                     := '0';             --       .oct_rzqin
		reset_reset_n      : in    std_logic                     := '0'              --  reset.reset_n
	);
end entity hps;

architecture rtl of hps is
	component hps_CNT_N is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component hps_CNT_N;

	component hps_K is
		port (
			clk         : in  std_logic                      := 'X';             -- clk
			address     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- address
			clken       : in  std_logic                      := 'X';             -- clken
			chipselect  : in  std_logic                      := 'X';             -- chipselect
			write       : in  std_logic                      := 'X';             -- write
			readdata    : out std_logic_vector(127 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                      := 'X';             -- reset
			reset_req   : in  std_logic                      := 'X';             -- reset_req
			address2    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- address
			chipselect2 : in  std_logic                      := 'X';             -- chipselect
			clken2      : in  std_logic                      := 'X';             -- clken
			write2      : in  std_logic                      := 'X';             -- write
			readdata2   : out std_logic_vector(127 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                      := 'X';             -- clk
			reset2      : in  std_logic                      := 'X';             -- reset
			reset_req2  : in  std_logic                      := 'X';             -- reset_req
			freeze      : in  std_logic                      := 'X'              -- freeze
		);
	end component hps_K;

	component hps_M is
		port (
			clk         : in  std_logic                      := 'X';             -- clk
			address     : in  std_logic_vector(9 downto 0)   := (others => 'X'); -- address
			clken       : in  std_logic                      := 'X';             -- clken
			chipselect  : in  std_logic                      := 'X';             -- chipselect
			write       : in  std_logic                      := 'X';             -- write
			readdata    : out std_logic_vector(127 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                      := 'X';             -- reset
			reset_req   : in  std_logic                      := 'X';             -- reset_req
			address2    : in  std_logic_vector(9 downto 0)   := (others => 'X'); -- address
			chipselect2 : in  std_logic                      := 'X';             -- chipselect
			clken2      : in  std_logic                      := 'X';             -- clken
			write2      : in  std_logic                      := 'X';             -- write
			readdata2   : out std_logic_vector(127 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                      := 'X';             -- clk
			reset2      : in  std_logic                      := 'X';             -- reset
			reset_req2  : in  std_logic                      := 'X';             -- reset_req
			freeze      : in  std_logic                      := 'X'              -- freeze
		);
	end component hps_M;

	component hps_a is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component hps_a;

	component hps_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			h2f_mpu_eventi     : in    std_logic                      := 'X';             -- eventi
			h2f_mpu_evento     : out   std_logic;                                         -- evento
			h2f_mpu_standbywfe : out   std_logic_vector(1 downto 0);                      -- standbywfe
			h2f_mpu_standbywfi : out   std_logic_vector(1 downto 0);                      -- standbywfi
			mem_a              : out   std_logic_vector(12 downto 0);                     -- mem_a
			mem_ba             : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck             : out   std_logic;                                         -- mem_ck
			mem_ck_n           : out   std_logic;                                         -- mem_ck_n
			mem_cke            : out   std_logic;                                         -- mem_cke
			mem_cs_n           : out   std_logic;                                         -- mem_cs_n
			mem_ras_n          : out   std_logic;                                         -- mem_ras_n
			mem_cas_n          : out   std_logic;                                         -- mem_cas_n
			mem_we_n           : out   std_logic;                                         -- mem_we_n
			mem_reset_n        : out   std_logic;                                         -- mem_reset_n
			mem_dq             : inout std_logic_vector(7 downto 0)   := (others => 'X'); -- mem_dq
			mem_dqs            : inout std_logic                      := 'X';             -- mem_dqs
			mem_dqs_n          : inout std_logic                      := 'X';             -- mem_dqs_n
			mem_odt            : out   std_logic;                                         -- mem_odt
			mem_dm             : out   std_logic;                                         -- mem_dm
			oct_rzqin          : in    std_logic                      := 'X';             -- oct_rzqin
			h2f_rst_n          : out   std_logic;                                         -- reset_n
			h2f_axi_clk        : in    std_logic                      := 'X';             -- clk
			h2f_AWID           : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR         : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN          : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE         : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST        : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK         : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE        : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT         : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID        : out   std_logic;                                         -- awvalid
			h2f_AWREADY        : in    std_logic                      := 'X';             -- awready
			h2f_WID            : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA          : out   std_logic_vector(127 downto 0);                    -- wdata
			h2f_WSTRB          : out   std_logic_vector(15 downto 0);                     -- wstrb
			h2f_WLAST          : out   std_logic;                                         -- wlast
			h2f_WVALID         : out   std_logic;                                         -- wvalid
			h2f_WREADY         : in    std_logic                      := 'X';             -- wready
			h2f_BID            : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP          : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID         : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY         : out   std_logic;                                         -- bready
			h2f_ARID           : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR         : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN          : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE         : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST        : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK         : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE        : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT         : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID        : out   std_logic;                                         -- arvalid
			h2f_ARREADY        : in    std_logic                      := 'X';             -- arready
			h2f_RID            : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA          : in    std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP          : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST          : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID         : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY         : out   std_logic;                                         -- rready
			h2f_lw_axi_clk     : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID        : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR      : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN       : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE      : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST     : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK      : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE     : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT      : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID     : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY     : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID         : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA       : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB       : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST       : out   std_logic;                                         -- wlast
			h2f_lw_WVALID      : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY      : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID         : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP       : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID      : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY      : out   std_logic;                                         -- bready
			h2f_lw_ARID        : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR      : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN       : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE      : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST     : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK      : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE     : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT      : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID     : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY     : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID         : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA       : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP       : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST       : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID      : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY      : out   std_logic;                                         -- rready
			f2h_irq_p0         : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- irq
			f2h_irq_p1         : in    std_logic_vector(31 downto 0)  := (others => 'X')  -- irq
		);
	end component hps_hps_0;

	component hps_interrupt is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			out_port   : out std_logic;                                        -- export
			irq        : out std_logic                                         -- irq
		);
	end component hps_interrupt;

	component hps_start is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			out_port   : out std_logic                                         -- export
		);
	end component hps_start;

	component hps_mm_interconnect_0 is
		port (
			hps_0_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- awid
			hps_0_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- awaddr
			hps_0_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			hps_0_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			hps_0_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			hps_0_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			hps_0_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			hps_0_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			hps_0_h2f_axi_master_awvalid                                     : in  std_logic                      := 'X';             -- awvalid
			hps_0_h2f_axi_master_awready                                     : out std_logic;                                         -- awready
			hps_0_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- wid
			hps_0_h2f_axi_master_wdata                                       : in  std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_axi_master_wstrb                                       : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_axi_master_wlast                                       : in  std_logic                      := 'X';             -- wlast
			hps_0_h2f_axi_master_wvalid                                      : in  std_logic                      := 'X';             -- wvalid
			hps_0_h2f_axi_master_wready                                      : out std_logic;                                         -- wready
			hps_0_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                     -- bid
			hps_0_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                      -- bresp
			hps_0_h2f_axi_master_bvalid                                      : out std_logic;                                         -- bvalid
			hps_0_h2f_axi_master_bready                                      : in  std_logic                      := 'X';             -- bready
			hps_0_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- arid
			hps_0_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- araddr
			hps_0_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			hps_0_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			hps_0_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			hps_0_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			hps_0_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			hps_0_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			hps_0_h2f_axi_master_arvalid                                     : in  std_logic                      := 'X';             -- arvalid
			hps_0_h2f_axi_master_arready                                     : out std_logic;                                         -- arready
			hps_0_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                     -- rid
			hps_0_h2f_axi_master_rdata                                       : out std_logic_vector(127 downto 0);                    -- rdata
			hps_0_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                      -- rresp
			hps_0_h2f_axi_master_rlast                                       : out std_logic;                                         -- rlast
			hps_0_h2f_axi_master_rvalid                                      : out std_logic;                                         -- rvalid
			hps_0_h2f_axi_master_rready                                      : in  std_logic                      := 'X';             -- rready
			clk_0_clk_clk                                                    : in  std_logic                      := 'X';             -- clk
			hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			K_reset1_reset_bridge_in_reset_reset                             : in  std_logic                      := 'X';             -- reset
			K_s1_address                                                     : out std_logic_vector(3 downto 0);                      -- address
			K_s1_write                                                       : out std_logic;                                         -- write
			K_s1_readdata                                                    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			K_s1_writedata                                                   : out std_logic_vector(127 downto 0);                    -- writedata
			K_s1_byteenable                                                  : out std_logic_vector(15 downto 0);                     -- byteenable
			K_s1_chipselect                                                  : out std_logic;                                         -- chipselect
			K_s1_clken                                                       : out std_logic;                                         -- clken
			M_s1_address                                                     : out std_logic_vector(9 downto 0);                      -- address
			M_s1_write                                                       : out std_logic;                                         -- write
			M_s1_readdata                                                    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			M_s1_writedata                                                   : out std_logic_vector(127 downto 0);                    -- writedata
			M_s1_byteenable                                                  : out std_logic_vector(15 downto 0);                     -- byteenable
			M_s1_chipselect                                                  : out std_logic;                                         -- chipselect
			M_s1_clken                                                       : out std_logic                                          -- clken
		);
	end component hps_mm_interconnect_0;

	component hps_mm_interconnect_1 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			CNT_N_reset_reset_bridge_in_reset_reset                             : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			a_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			a_s1_write                                                          : out std_logic;                                        -- write
			a_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			a_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			a_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			a_init_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			a_init_s1_write                                                     : out std_logic;                                        -- write
			a_init_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			a_init_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			a_init_s1_chipselect                                                : out std_logic;                                        -- chipselect
			b_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			b_s1_write                                                          : out std_logic;                                        -- write
			b_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			b_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			b_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			b_init_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			b_init_s1_write                                                     : out std_logic;                                        -- write
			b_init_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			b_init_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			b_init_s1_chipselect                                                : out std_logic;                                        -- chipselect
			c_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			c_s1_write                                                          : out std_logic;                                        -- write
			c_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			c_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			c_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			c_init_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			c_init_s1_write                                                     : out std_logic;                                        -- write
			c_init_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			c_init_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			c_init_s1_chipselect                                                : out std_logic;                                        -- chipselect
			CNT_N_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			CNT_N_s1_write                                                      : out std_logic;                                        -- write
			CNT_N_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CNT_N_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			CNT_N_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			d_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			d_s1_write                                                          : out std_logic;                                        -- write
			d_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			d_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			d_init_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			d_init_s1_write                                                     : out std_logic;                                        -- write
			d_init_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_init_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			d_init_s1_chipselect                                                : out std_logic;                                        -- chipselect
			e_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			e_s1_write                                                          : out std_logic;                                        -- write
			e_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			e_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			e_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			e_init_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			e_init_s1_write                                                     : out std_logic;                                        -- write
			e_init_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			e_init_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			e_init_s1_chipselect                                                : out std_logic;                                        -- chipselect
			f_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			f_s1_write                                                          : out std_logic;                                        -- write
			f_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			f_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			f_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			f_init_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			f_init_s1_write                                                     : out std_logic;                                        -- write
			f_init_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			f_init_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			f_init_s1_chipselect                                                : out std_logic;                                        -- chipselect
			g_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			g_s1_write                                                          : out std_logic;                                        -- write
			g_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			g_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			g_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			g_init_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			g_init_s1_write                                                     : out std_logic;                                        -- write
			g_init_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			g_init_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			g_init_s1_chipselect                                                : out std_logic;                                        -- chipselect
			h_s1_address                                                        : out std_logic_vector(1 downto 0);                     -- address
			h_s1_write                                                          : out std_logic;                                        -- write
			h_s1_readdata                                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			h_s1_writedata                                                      : out std_logic_vector(31 downto 0);                    -- writedata
			h_s1_chipselect                                                     : out std_logic;                                        -- chipselect
			h_init_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			h_init_s1_write                                                     : out std_logic;                                        -- write
			h_init_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			h_init_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			h_init_s1_chipselect                                                : out std_logic;                                        -- chipselect
			interrupt_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			interrupt_s1_write                                                  : out std_logic;                                        -- write
			interrupt_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			interrupt_s1_writedata                                              : out std_logic_vector(31 downto 0);                    -- writedata
			interrupt_s1_chipselect                                             : out std_logic;                                        -- chipselect
			start_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			start_s1_write                                                      : out std_logic;                                        -- write
			start_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			start_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			start_s1_chipselect                                                 : out std_logic                                         -- chipselect
		);
	end component hps_mm_interconnect_1;

	component hps_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component hps_irq_mapper;

	component hps_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component hps_irq_mapper_001;

	component hps_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component hps_rst_controller;

	component hps_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component hps_rst_controller_001;

	signal hps_0_h2f_axi_master_awburst                   : std_logic_vector(1 downto 0);   -- hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	signal hps_0_h2f_axi_master_arlen                     : std_logic_vector(3 downto 0);   -- hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	signal hps_0_h2f_axi_master_wstrb                     : std_logic_vector(15 downto 0);  -- hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	signal hps_0_h2f_axi_master_wready                    : std_logic;                      -- mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	signal hps_0_h2f_axi_master_rid                       : std_logic_vector(11 downto 0);  -- mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	signal hps_0_h2f_axi_master_rready                    : std_logic;                      -- hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	signal hps_0_h2f_axi_master_awlen                     : std_logic_vector(3 downto 0);   -- hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	signal hps_0_h2f_axi_master_wid                       : std_logic_vector(11 downto 0);  -- hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	signal hps_0_h2f_axi_master_arcache                   : std_logic_vector(3 downto 0);   -- hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	signal hps_0_h2f_axi_master_wvalid                    : std_logic;                      -- hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	signal hps_0_h2f_axi_master_araddr                    : std_logic_vector(29 downto 0);  -- hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	signal hps_0_h2f_axi_master_arprot                    : std_logic_vector(2 downto 0);   -- hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	signal hps_0_h2f_axi_master_awprot                    : std_logic_vector(2 downto 0);   -- hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	signal hps_0_h2f_axi_master_wdata                     : std_logic_vector(127 downto 0); -- hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	signal hps_0_h2f_axi_master_arvalid                   : std_logic;                      -- hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	signal hps_0_h2f_axi_master_awcache                   : std_logic_vector(3 downto 0);   -- hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	signal hps_0_h2f_axi_master_arid                      : std_logic_vector(11 downto 0);  -- hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	signal hps_0_h2f_axi_master_arlock                    : std_logic_vector(1 downto 0);   -- hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	signal hps_0_h2f_axi_master_awlock                    : std_logic_vector(1 downto 0);   -- hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	signal hps_0_h2f_axi_master_awaddr                    : std_logic_vector(29 downto 0);  -- hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	signal hps_0_h2f_axi_master_bresp                     : std_logic_vector(1 downto 0);   -- mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	signal hps_0_h2f_axi_master_arready                   : std_logic;                      -- mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	signal hps_0_h2f_axi_master_rdata                     : std_logic_vector(127 downto 0); -- mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	signal hps_0_h2f_axi_master_awready                   : std_logic;                      -- mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	signal hps_0_h2f_axi_master_arburst                   : std_logic_vector(1 downto 0);   -- hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	signal hps_0_h2f_axi_master_arsize                    : std_logic_vector(2 downto 0);   -- hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	signal hps_0_h2f_axi_master_bready                    : std_logic;                      -- hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	signal hps_0_h2f_axi_master_rlast                     : std_logic;                      -- mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	signal hps_0_h2f_axi_master_wlast                     : std_logic;                      -- hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	signal hps_0_h2f_axi_master_rresp                     : std_logic_vector(1 downto 0);   -- mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	signal hps_0_h2f_axi_master_awid                      : std_logic_vector(11 downto 0);  -- hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	signal hps_0_h2f_axi_master_bid                       : std_logic_vector(11 downto 0);  -- mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	signal hps_0_h2f_axi_master_bvalid                    : std_logic;                      -- mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	signal hps_0_h2f_axi_master_awsize                    : std_logic_vector(2 downto 0);   -- hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	signal hps_0_h2f_axi_master_awvalid                   : std_logic;                      -- hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	signal hps_0_h2f_axi_master_rvalid                    : std_logic;                      -- mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	signal mm_interconnect_0_k_s1_chipselect              : std_logic;                      -- mm_interconnect_0:K_s1_chipselect -> K:chipselect
	signal mm_interconnect_0_k_s1_readdata                : std_logic_vector(127 downto 0); -- K:readdata -> mm_interconnect_0:K_s1_readdata
	signal mm_interconnect_0_k_s1_address                 : std_logic_vector(3 downto 0);   -- mm_interconnect_0:K_s1_address -> K:address
	signal mm_interconnect_0_k_s1_byteenable              : std_logic_vector(15 downto 0);  -- mm_interconnect_0:K_s1_byteenable -> K:byteenable
	signal mm_interconnect_0_k_s1_write                   : std_logic;                      -- mm_interconnect_0:K_s1_write -> K:write
	signal mm_interconnect_0_k_s1_writedata               : std_logic_vector(127 downto 0); -- mm_interconnect_0:K_s1_writedata -> K:writedata
	signal mm_interconnect_0_k_s1_clken                   : std_logic;                      -- mm_interconnect_0:K_s1_clken -> K:clken
	signal mm_interconnect_0_m_s1_chipselect              : std_logic;                      -- mm_interconnect_0:M_s1_chipselect -> M:chipselect
	signal mm_interconnect_0_m_s1_readdata                : std_logic_vector(127 downto 0); -- M:readdata -> mm_interconnect_0:M_s1_readdata
	signal mm_interconnect_0_m_s1_address                 : std_logic_vector(9 downto 0);   -- mm_interconnect_0:M_s1_address -> M:address
	signal mm_interconnect_0_m_s1_byteenable              : std_logic_vector(15 downto 0);  -- mm_interconnect_0:M_s1_byteenable -> M:byteenable
	signal mm_interconnect_0_m_s1_write                   : std_logic;                      -- mm_interconnect_0:M_s1_write -> M:write
	signal mm_interconnect_0_m_s1_writedata               : std_logic_vector(127 downto 0); -- mm_interconnect_0:M_s1_writedata -> M:writedata
	signal mm_interconnect_0_m_s1_clken                   : std_logic;                      -- mm_interconnect_0:M_s1_clken -> M:clken
	signal hps_0_h2f_lw_axi_master_awburst                : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                  : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                  : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                 : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                    : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                 : std_logic;                      -- hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                  : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                    : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                 : std_logic;                      -- hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                 : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                 : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                 : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                  : std_logic_vector(31 downto 0);  -- hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                : std_logic;                      -- hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                   : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                 : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                 : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                 : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                  : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                  : std_logic_vector(31 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                 : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                 : std_logic;                      -- hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                  : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                  : std_logic;                      -- hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                  : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                   : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                    : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                 : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                 : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                : std_logic;                      -- hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                 : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_1_cnt_n_s1_chipselect          : std_logic;                      -- mm_interconnect_1:CNT_N_s1_chipselect -> CNT_N:chipselect
	signal mm_interconnect_1_cnt_n_s1_readdata            : std_logic_vector(31 downto 0);  -- CNT_N:readdata -> mm_interconnect_1:CNT_N_s1_readdata
	signal mm_interconnect_1_cnt_n_s1_address             : std_logic_vector(1 downto 0);   -- mm_interconnect_1:CNT_N_s1_address -> CNT_N:address
	signal mm_interconnect_1_cnt_n_s1_write               : std_logic;                      -- mm_interconnect_1:CNT_N_s1_write -> mm_interconnect_1_cnt_n_s1_write:in
	signal mm_interconnect_1_cnt_n_s1_writedata           : std_logic_vector(31 downto 0);  -- mm_interconnect_1:CNT_N_s1_writedata -> CNT_N:writedata
	signal mm_interconnect_1_a_init_s1_chipselect         : std_logic;                      -- mm_interconnect_1:a_init_s1_chipselect -> a_init:chipselect
	signal mm_interconnect_1_a_init_s1_readdata           : std_logic_vector(31 downto 0);  -- a_init:readdata -> mm_interconnect_1:a_init_s1_readdata
	signal mm_interconnect_1_a_init_s1_address            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:a_init_s1_address -> a_init:address
	signal mm_interconnect_1_a_init_s1_write              : std_logic;                      -- mm_interconnect_1:a_init_s1_write -> mm_interconnect_1_a_init_s1_write:in
	signal mm_interconnect_1_a_init_s1_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:a_init_s1_writedata -> a_init:writedata
	signal mm_interconnect_1_b_init_s1_chipselect         : std_logic;                      -- mm_interconnect_1:b_init_s1_chipselect -> b_init:chipselect
	signal mm_interconnect_1_b_init_s1_readdata           : std_logic_vector(31 downto 0);  -- b_init:readdata -> mm_interconnect_1:b_init_s1_readdata
	signal mm_interconnect_1_b_init_s1_address            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:b_init_s1_address -> b_init:address
	signal mm_interconnect_1_b_init_s1_write              : std_logic;                      -- mm_interconnect_1:b_init_s1_write -> mm_interconnect_1_b_init_s1_write:in
	signal mm_interconnect_1_b_init_s1_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:b_init_s1_writedata -> b_init:writedata
	signal mm_interconnect_1_c_init_s1_chipselect         : std_logic;                      -- mm_interconnect_1:c_init_s1_chipselect -> c_init:chipselect
	signal mm_interconnect_1_c_init_s1_readdata           : std_logic_vector(31 downto 0);  -- c_init:readdata -> mm_interconnect_1:c_init_s1_readdata
	signal mm_interconnect_1_c_init_s1_address            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:c_init_s1_address -> c_init:address
	signal mm_interconnect_1_c_init_s1_write              : std_logic;                      -- mm_interconnect_1:c_init_s1_write -> mm_interconnect_1_c_init_s1_write:in
	signal mm_interconnect_1_c_init_s1_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:c_init_s1_writedata -> c_init:writedata
	signal mm_interconnect_1_d_init_s1_chipselect         : std_logic;                      -- mm_interconnect_1:d_init_s1_chipselect -> d_init:chipselect
	signal mm_interconnect_1_d_init_s1_readdata           : std_logic_vector(31 downto 0);  -- d_init:readdata -> mm_interconnect_1:d_init_s1_readdata
	signal mm_interconnect_1_d_init_s1_address            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:d_init_s1_address -> d_init:address
	signal mm_interconnect_1_d_init_s1_write              : std_logic;                      -- mm_interconnect_1:d_init_s1_write -> mm_interconnect_1_d_init_s1_write:in
	signal mm_interconnect_1_d_init_s1_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:d_init_s1_writedata -> d_init:writedata
	signal mm_interconnect_1_e_init_s1_chipselect         : std_logic;                      -- mm_interconnect_1:e_init_s1_chipselect -> e_init:chipselect
	signal mm_interconnect_1_e_init_s1_readdata           : std_logic_vector(31 downto 0);  -- e_init:readdata -> mm_interconnect_1:e_init_s1_readdata
	signal mm_interconnect_1_e_init_s1_address            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:e_init_s1_address -> e_init:address
	signal mm_interconnect_1_e_init_s1_write              : std_logic;                      -- mm_interconnect_1:e_init_s1_write -> mm_interconnect_1_e_init_s1_write:in
	signal mm_interconnect_1_e_init_s1_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:e_init_s1_writedata -> e_init:writedata
	signal mm_interconnect_1_f_init_s1_chipselect         : std_logic;                      -- mm_interconnect_1:f_init_s1_chipselect -> f_init:chipselect
	signal mm_interconnect_1_f_init_s1_readdata           : std_logic_vector(31 downto 0);  -- f_init:readdata -> mm_interconnect_1:f_init_s1_readdata
	signal mm_interconnect_1_f_init_s1_address            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:f_init_s1_address -> f_init:address
	signal mm_interconnect_1_f_init_s1_write              : std_logic;                      -- mm_interconnect_1:f_init_s1_write -> mm_interconnect_1_f_init_s1_write:in
	signal mm_interconnect_1_f_init_s1_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:f_init_s1_writedata -> f_init:writedata
	signal mm_interconnect_1_g_init_s1_chipselect         : std_logic;                      -- mm_interconnect_1:g_init_s1_chipselect -> g_init:chipselect
	signal mm_interconnect_1_g_init_s1_readdata           : std_logic_vector(31 downto 0);  -- g_init:readdata -> mm_interconnect_1:g_init_s1_readdata
	signal mm_interconnect_1_g_init_s1_address            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:g_init_s1_address -> g_init:address
	signal mm_interconnect_1_g_init_s1_write              : std_logic;                      -- mm_interconnect_1:g_init_s1_write -> mm_interconnect_1_g_init_s1_write:in
	signal mm_interconnect_1_g_init_s1_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:g_init_s1_writedata -> g_init:writedata
	signal mm_interconnect_1_h_init_s1_chipselect         : std_logic;                      -- mm_interconnect_1:h_init_s1_chipselect -> h_init:chipselect
	signal mm_interconnect_1_h_init_s1_readdata           : std_logic_vector(31 downto 0);  -- h_init:readdata -> mm_interconnect_1:h_init_s1_readdata
	signal mm_interconnect_1_h_init_s1_address            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:h_init_s1_address -> h_init:address
	signal mm_interconnect_1_h_init_s1_write              : std_logic;                      -- mm_interconnect_1:h_init_s1_write -> mm_interconnect_1_h_init_s1_write:in
	signal mm_interconnect_1_h_init_s1_writedata          : std_logic_vector(31 downto 0);  -- mm_interconnect_1:h_init_s1_writedata -> h_init:writedata
	signal mm_interconnect_1_a_s1_chipselect              : std_logic;                      -- mm_interconnect_1:a_s1_chipselect -> a:chipselect
	signal mm_interconnect_1_a_s1_readdata                : std_logic_vector(31 downto 0);  -- a:readdata -> mm_interconnect_1:a_s1_readdata
	signal mm_interconnect_1_a_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:a_s1_address -> a:address
	signal mm_interconnect_1_a_s1_write                   : std_logic;                      -- mm_interconnect_1:a_s1_write -> mm_interconnect_1_a_s1_write:in
	signal mm_interconnect_1_a_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:a_s1_writedata -> a:writedata
	signal mm_interconnect_1_b_s1_chipselect              : std_logic;                      -- mm_interconnect_1:b_s1_chipselect -> b:chipselect
	signal mm_interconnect_1_b_s1_readdata                : std_logic_vector(31 downto 0);  -- b:readdata -> mm_interconnect_1:b_s1_readdata
	signal mm_interconnect_1_b_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:b_s1_address -> b:address
	signal mm_interconnect_1_b_s1_write                   : std_logic;                      -- mm_interconnect_1:b_s1_write -> mm_interconnect_1_b_s1_write:in
	signal mm_interconnect_1_b_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:b_s1_writedata -> b:writedata
	signal mm_interconnect_1_c_s1_chipselect              : std_logic;                      -- mm_interconnect_1:c_s1_chipselect -> c:chipselect
	signal mm_interconnect_1_c_s1_readdata                : std_logic_vector(31 downto 0);  -- c:readdata -> mm_interconnect_1:c_s1_readdata
	signal mm_interconnect_1_c_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:c_s1_address -> c:address
	signal mm_interconnect_1_c_s1_write                   : std_logic;                      -- mm_interconnect_1:c_s1_write -> mm_interconnect_1_c_s1_write:in
	signal mm_interconnect_1_c_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:c_s1_writedata -> c:writedata
	signal mm_interconnect_1_d_s1_chipselect              : std_logic;                      -- mm_interconnect_1:d_s1_chipselect -> d:chipselect
	signal mm_interconnect_1_d_s1_readdata                : std_logic_vector(31 downto 0);  -- d:readdata -> mm_interconnect_1:d_s1_readdata
	signal mm_interconnect_1_d_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:d_s1_address -> d:address
	signal mm_interconnect_1_d_s1_write                   : std_logic;                      -- mm_interconnect_1:d_s1_write -> mm_interconnect_1_d_s1_write:in
	signal mm_interconnect_1_d_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:d_s1_writedata -> d:writedata
	signal mm_interconnect_1_e_s1_chipselect              : std_logic;                      -- mm_interconnect_1:e_s1_chipselect -> e:chipselect
	signal mm_interconnect_1_e_s1_readdata                : std_logic_vector(31 downto 0);  -- e:readdata -> mm_interconnect_1:e_s1_readdata
	signal mm_interconnect_1_e_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:e_s1_address -> e:address
	signal mm_interconnect_1_e_s1_write                   : std_logic;                      -- mm_interconnect_1:e_s1_write -> mm_interconnect_1_e_s1_write:in
	signal mm_interconnect_1_e_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:e_s1_writedata -> e:writedata
	signal mm_interconnect_1_f_s1_chipselect              : std_logic;                      -- mm_interconnect_1:f_s1_chipselect -> f:chipselect
	signal mm_interconnect_1_f_s1_readdata                : std_logic_vector(31 downto 0);  -- f:readdata -> mm_interconnect_1:f_s1_readdata
	signal mm_interconnect_1_f_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:f_s1_address -> f:address
	signal mm_interconnect_1_f_s1_write                   : std_logic;                      -- mm_interconnect_1:f_s1_write -> mm_interconnect_1_f_s1_write:in
	signal mm_interconnect_1_f_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:f_s1_writedata -> f:writedata
	signal mm_interconnect_1_g_s1_chipselect              : std_logic;                      -- mm_interconnect_1:g_s1_chipselect -> g:chipselect
	signal mm_interconnect_1_g_s1_readdata                : std_logic_vector(31 downto 0);  -- g:readdata -> mm_interconnect_1:g_s1_readdata
	signal mm_interconnect_1_g_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:g_s1_address -> g:address
	signal mm_interconnect_1_g_s1_write                   : std_logic;                      -- mm_interconnect_1:g_s1_write -> mm_interconnect_1_g_s1_write:in
	signal mm_interconnect_1_g_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:g_s1_writedata -> g:writedata
	signal mm_interconnect_1_h_s1_chipselect              : std_logic;                      -- mm_interconnect_1:h_s1_chipselect -> h:chipselect
	signal mm_interconnect_1_h_s1_readdata                : std_logic_vector(31 downto 0);  -- h:readdata -> mm_interconnect_1:h_s1_readdata
	signal mm_interconnect_1_h_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:h_s1_address -> h:address
	signal mm_interconnect_1_h_s1_write                   : std_logic;                      -- mm_interconnect_1:h_s1_write -> mm_interconnect_1_h_s1_write:in
	signal mm_interconnect_1_h_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:h_s1_writedata -> h:writedata
	signal mm_interconnect_1_start_s1_chipselect          : std_logic;                      -- mm_interconnect_1:start_s1_chipselect -> start:chipselect
	signal mm_interconnect_1_start_s1_readdata            : std_logic_vector(31 downto 0);  -- start:readdata -> mm_interconnect_1:start_s1_readdata
	signal mm_interconnect_1_start_s1_address             : std_logic_vector(1 downto 0);   -- mm_interconnect_1:start_s1_address -> start:address
	signal mm_interconnect_1_start_s1_write               : std_logic;                      -- mm_interconnect_1:start_s1_write -> mm_interconnect_1_start_s1_write:in
	signal mm_interconnect_1_start_s1_writedata           : std_logic_vector(31 downto 0);  -- mm_interconnect_1:start_s1_writedata -> start:writedata
	signal mm_interconnect_1_interrupt_s1_chipselect      : std_logic;                      -- mm_interconnect_1:interrupt_s1_chipselect -> interrupt:chipselect
	signal mm_interconnect_1_interrupt_s1_readdata        : std_logic_vector(31 downto 0);  -- interrupt:readdata -> mm_interconnect_1:interrupt_s1_readdata
	signal mm_interconnect_1_interrupt_s1_address         : std_logic_vector(1 downto 0);   -- mm_interconnect_1:interrupt_s1_address -> interrupt:address
	signal mm_interconnect_1_interrupt_s1_write           : std_logic;                      -- mm_interconnect_1:interrupt_s1_write -> mm_interconnect_1_interrupt_s1_write:in
	signal mm_interconnect_1_interrupt_s1_writedata       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:interrupt_s1_writedata -> interrupt:writedata
	signal irq_mapper_receiver0_irq                       : std_logic;                      -- interrupt:irq -> irq_mapper:receiver0_irq
	signal hps_0_f2h_irq0_irq                             : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	signal hps_0_f2h_irq1_irq                             : std_logic_vector(31 downto 0);  -- irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	signal rst_controller_reset_out_reset                 : std_logic;                      -- rst_controller:reset_out -> [K:reset, K:reset2, M:reset, M:reset2, mm_interconnect_0:K_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:CNT_N_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req             : std_logic;                      -- rst_controller:reset_req -> [K:reset_req, K:reset_req2, M:reset_req, M:reset_req2, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset             : std_logic;                      -- rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal hps_0_h2f_reset_reset                          : std_logic;                      -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal reset_reset_n_ports_inv                        : std_logic;                      -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_1_cnt_n_s1_write_ports_inv     : std_logic;                      -- mm_interconnect_1_cnt_n_s1_write:inv -> CNT_N:write_n
	signal mm_interconnect_1_a_init_s1_write_ports_inv    : std_logic;                      -- mm_interconnect_1_a_init_s1_write:inv -> a_init:write_n
	signal mm_interconnect_1_b_init_s1_write_ports_inv    : std_logic;                      -- mm_interconnect_1_b_init_s1_write:inv -> b_init:write_n
	signal mm_interconnect_1_c_init_s1_write_ports_inv    : std_logic;                      -- mm_interconnect_1_c_init_s1_write:inv -> c_init:write_n
	signal mm_interconnect_1_d_init_s1_write_ports_inv    : std_logic;                      -- mm_interconnect_1_d_init_s1_write:inv -> d_init:write_n
	signal mm_interconnect_1_e_init_s1_write_ports_inv    : std_logic;                      -- mm_interconnect_1_e_init_s1_write:inv -> e_init:write_n
	signal mm_interconnect_1_f_init_s1_write_ports_inv    : std_logic;                      -- mm_interconnect_1_f_init_s1_write:inv -> f_init:write_n
	signal mm_interconnect_1_g_init_s1_write_ports_inv    : std_logic;                      -- mm_interconnect_1_g_init_s1_write:inv -> g_init:write_n
	signal mm_interconnect_1_h_init_s1_write_ports_inv    : std_logic;                      -- mm_interconnect_1_h_init_s1_write:inv -> h_init:write_n
	signal mm_interconnect_1_a_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_a_s1_write:inv -> a:write_n
	signal mm_interconnect_1_b_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_b_s1_write:inv -> b:write_n
	signal mm_interconnect_1_c_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_c_s1_write:inv -> c:write_n
	signal mm_interconnect_1_d_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_d_s1_write:inv -> d:write_n
	signal mm_interconnect_1_e_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_e_s1_write:inv -> e:write_n
	signal mm_interconnect_1_f_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_f_s1_write:inv -> f:write_n
	signal mm_interconnect_1_g_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_g_s1_write:inv -> g:write_n
	signal mm_interconnect_1_h_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_h_s1_write:inv -> h:write_n
	signal mm_interconnect_1_start_s1_write_ports_inv     : std_logic;                      -- mm_interconnect_1_start_s1_write:inv -> start:write_n
	signal mm_interconnect_1_interrupt_s1_write_ports_inv : std_logic;                      -- mm_interconnect_1_interrupt_s1_write:inv -> interrupt:write_n
	signal rst_controller_reset_out_reset_ports_inv       : std_logic;                      -- rst_controller_reset_out_reset:inv -> [CNT_N:reset_n, a:reset_n, a_init:reset_n, b:reset_n, b_init:reset_n, c:reset_n, c_init:reset_n, d:reset_n, d_init:reset_n, e:reset_n, e_init:reset_n, f:reset_n, f_init:reset_n, g:reset_n, g_init:reset_n, h:reset_n, h_init:reset_n, interrupt:reset_n, start:reset_n]
	signal hps_0_h2f_reset_reset_ports_inv                : std_logic;                      -- hps_0_h2f_reset_reset:inv -> rst_controller_001:reset_in0

begin

	cnt_n : component hps_CNT_N
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_1_cnt_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_cnt_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_cnt_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_cnt_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_cnt_n_s1_readdata,        --                    .readdata
			in_port    => open,                                       -- external_connection.export
			out_port   => open                                        --                    .export
		);

	k : component hps_K
		port map (
			clk         => clk_clk,                            --   clk1.clk
			address     => mm_interconnect_0_k_s1_address,     --     s1.address
			clken       => mm_interconnect_0_k_s1_clken,       --       .clken
			chipselect  => mm_interconnect_0_k_s1_chipselect,  --       .chipselect
			write       => mm_interconnect_0_k_s1_write,       --       .write
			readdata    => mm_interconnect_0_k_s1_readdata,    --       .readdata
			writedata   => mm_interconnect_0_k_s1_writedata,   --       .writedata
			byteenable  => mm_interconnect_0_k_s1_byteenable,  --       .byteenable
			reset       => rst_controller_reset_out_reset,     -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req, --       .reset_req
			address2    => open,                               --     s2.address
			chipselect2 => open,                               --       .chipselect
			clken2      => open,                               --       .clken
			write2      => open,                               --       .write
			readdata2   => open,                               --       .readdata
			writedata2  => open,                               --       .writedata
			byteenable2 => open,                               --       .byteenable
			clk2        => clk_clk,                            --   clk2.clk
			reset2      => rst_controller_reset_out_reset,     -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req, --       .reset_req
			freeze      => '0'                                 -- (terminated)
		);

	m : component hps_M
		port map (
			clk         => clk_clk,                            --   clk1.clk
			address     => mm_interconnect_0_m_s1_address,     --     s1.address
			clken       => mm_interconnect_0_m_s1_clken,       --       .clken
			chipselect  => mm_interconnect_0_m_s1_chipselect,  --       .chipselect
			write       => mm_interconnect_0_m_s1_write,       --       .write
			readdata    => mm_interconnect_0_m_s1_readdata,    --       .readdata
			writedata   => mm_interconnect_0_m_s1_writedata,   --       .writedata
			byteenable  => mm_interconnect_0_m_s1_byteenable,  --       .byteenable
			reset       => rst_controller_reset_out_reset,     -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req, --       .reset_req
			address2    => open,                               --     s2.address
			chipselect2 => open,                               --       .chipselect
			clken2      => open,                               --       .clken
			write2      => open,                               --       .write
			readdata2   => open,                               --       .readdata
			writedata2  => open,                               --       .writedata
			byteenable2 => open,                               --       .byteenable
			clk2        => clk_clk,                            --   clk2.clk
			reset2      => rst_controller_reset_out_reset,     -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req, --       .reset_req
			freeze      => '0'                                 -- (terminated)
		);

	a : component hps_a
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_a_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_a_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_a_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_a_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_a_s1_readdata,          --                    .readdata
			in_port    => open,                                     -- external_connection.export
			out_port   => open                                      --                    .export
		);

	a_init : component hps_a
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_a_init_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_a_init_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_a_init_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_a_init_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_a_init_s1_readdata,        --                    .readdata
			in_port    => open,                                        -- external_connection.export
			out_port   => open                                         --                    .export
		);

	b : component hps_a
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_b_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_b_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_b_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_b_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_b_s1_readdata,          --                    .readdata
			in_port    => open,                                     -- external_connection.export
			out_port   => open                                      --                    .export
		);

	b_init : component hps_a
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_b_init_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_b_init_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_b_init_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_b_init_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_b_init_s1_readdata,        --                    .readdata
			in_port    => open,                                        -- external_connection.export
			out_port   => open                                         --                    .export
		);

	c : component hps_a
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_c_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_c_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_c_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_c_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_c_s1_readdata,          --                    .readdata
			in_port    => open,                                     -- external_connection.export
			out_port   => open                                      --                    .export
		);

	c_init : component hps_a
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_c_init_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_c_init_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_c_init_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_c_init_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_c_init_s1_readdata,        --                    .readdata
			in_port    => open,                                        -- external_connection.export
			out_port   => open                                         --                    .export
		);

	d : component hps_a
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_d_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_d_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_d_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_d_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_d_s1_readdata,          --                    .readdata
			in_port    => open,                                     -- external_connection.export
			out_port   => open                                      --                    .export
		);

	d_init : component hps_a
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_d_init_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_d_init_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_d_init_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_d_init_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_d_init_s1_readdata,        --                    .readdata
			in_port    => open,                                        -- external_connection.export
			out_port   => open                                         --                    .export
		);

	e : component hps_a
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_e_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_e_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_e_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_e_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_e_s1_readdata,          --                    .readdata
			in_port    => open,                                     -- external_connection.export
			out_port   => open                                      --                    .export
		);

	e_init : component hps_a
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_e_init_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_e_init_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_e_init_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_e_init_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_e_init_s1_readdata,        --                    .readdata
			in_port    => open,                                        -- external_connection.export
			out_port   => open                                         --                    .export
		);

	f : component hps_a
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_f_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_f_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_f_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_f_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_f_s1_readdata,          --                    .readdata
			in_port    => open,                                     -- external_connection.export
			out_port   => open                                      --                    .export
		);

	f_init : component hps_a
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_f_init_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_f_init_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_f_init_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_f_init_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_f_init_s1_readdata,        --                    .readdata
			in_port    => open,                                        -- external_connection.export
			out_port   => open                                         --                    .export
		);

	g : component hps_a
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_g_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_g_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_g_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_g_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_g_s1_readdata,          --                    .readdata
			in_port    => open,                                     -- external_connection.export
			out_port   => open                                      --                    .export
		);

	g_init : component hps_a
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_g_init_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_g_init_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_g_init_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_g_init_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_g_init_s1_readdata,        --                    .readdata
			in_port    => open,                                        -- external_connection.export
			out_port   => open                                         --                    .export
		);

	h : component hps_a
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_1_h_s1_address,           --                  s1.address
			write_n    => mm_interconnect_1_h_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_1_h_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_1_h_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_1_h_s1_readdata,          --                    .readdata
			in_port    => open,                                     -- external_connection.export
			out_port   => open                                      --                    .export
		);

	h_init : component hps_a
		port map (
			clk        => clk_clk,                                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_1_h_init_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_h_init_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_h_init_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_h_init_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_h_init_s1_readdata,        --                    .readdata
			in_port    => open,                                        -- external_connection.export
			out_port   => open                                         --                    .export
		);

	hps_0 : component hps_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 3
		)
		port map (
			h2f_mpu_eventi     => open,                            --    h2f_mpu_events.eventi
			h2f_mpu_evento     => open,                            --                  .evento
			h2f_mpu_standbywfe => open,                            --                  .standbywfe
			h2f_mpu_standbywfi => open,                            --                  .standbywfi
			mem_a              => memory_mem_a,                    --            memory.mem_a
			mem_ba             => memory_mem_ba,                   --                  .mem_ba
			mem_ck             => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n           => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke            => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n           => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n          => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n          => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n           => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n        => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq             => memory_mem_dq,                   --                  .mem_dq
			mem_dqs            => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n          => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt            => memory_mem_odt,                  --                  .mem_odt
			mem_dm             => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin          => memory_oct_rzqin,                --                  .oct_rzqin
			h2f_rst_n          => hps_0_h2f_reset_reset,           --         h2f_reset.reset_n
			h2f_axi_clk        => clk_clk,                         --     h2f_axi_clock.clk
			h2f_AWID           => hps_0_h2f_axi_master_awid,       --    h2f_axi_master.awid
			h2f_AWADDR         => hps_0_h2f_axi_master_awaddr,     --                  .awaddr
			h2f_AWLEN          => hps_0_h2f_axi_master_awlen,      --                  .awlen
			h2f_AWSIZE         => hps_0_h2f_axi_master_awsize,     --                  .awsize
			h2f_AWBURST        => hps_0_h2f_axi_master_awburst,    --                  .awburst
			h2f_AWLOCK         => hps_0_h2f_axi_master_awlock,     --                  .awlock
			h2f_AWCACHE        => hps_0_h2f_axi_master_awcache,    --                  .awcache
			h2f_AWPROT         => hps_0_h2f_axi_master_awprot,     --                  .awprot
			h2f_AWVALID        => hps_0_h2f_axi_master_awvalid,    --                  .awvalid
			h2f_AWREADY        => hps_0_h2f_axi_master_awready,    --                  .awready
			h2f_WID            => hps_0_h2f_axi_master_wid,        --                  .wid
			h2f_WDATA          => hps_0_h2f_axi_master_wdata,      --                  .wdata
			h2f_WSTRB          => hps_0_h2f_axi_master_wstrb,      --                  .wstrb
			h2f_WLAST          => hps_0_h2f_axi_master_wlast,      --                  .wlast
			h2f_WVALID         => hps_0_h2f_axi_master_wvalid,     --                  .wvalid
			h2f_WREADY         => hps_0_h2f_axi_master_wready,     --                  .wready
			h2f_BID            => hps_0_h2f_axi_master_bid,        --                  .bid
			h2f_BRESP          => hps_0_h2f_axi_master_bresp,      --                  .bresp
			h2f_BVALID         => hps_0_h2f_axi_master_bvalid,     --                  .bvalid
			h2f_BREADY         => hps_0_h2f_axi_master_bready,     --                  .bready
			h2f_ARID           => hps_0_h2f_axi_master_arid,       --                  .arid
			h2f_ARADDR         => hps_0_h2f_axi_master_araddr,     --                  .araddr
			h2f_ARLEN          => hps_0_h2f_axi_master_arlen,      --                  .arlen
			h2f_ARSIZE         => hps_0_h2f_axi_master_arsize,     --                  .arsize
			h2f_ARBURST        => hps_0_h2f_axi_master_arburst,    --                  .arburst
			h2f_ARLOCK         => hps_0_h2f_axi_master_arlock,     --                  .arlock
			h2f_ARCACHE        => hps_0_h2f_axi_master_arcache,    --                  .arcache
			h2f_ARPROT         => hps_0_h2f_axi_master_arprot,     --                  .arprot
			h2f_ARVALID        => hps_0_h2f_axi_master_arvalid,    --                  .arvalid
			h2f_ARREADY        => hps_0_h2f_axi_master_arready,    --                  .arready
			h2f_RID            => hps_0_h2f_axi_master_rid,        --                  .rid
			h2f_RDATA          => hps_0_h2f_axi_master_rdata,      --                  .rdata
			h2f_RRESP          => hps_0_h2f_axi_master_rresp,      --                  .rresp
			h2f_RLAST          => hps_0_h2f_axi_master_rlast,      --                  .rlast
			h2f_RVALID         => hps_0_h2f_axi_master_rvalid,     --                  .rvalid
			h2f_RREADY         => hps_0_h2f_axi_master_rready,     --                  .rready
			h2f_lw_axi_clk     => clk_clk,                         --  h2f_lw_axi_clock.clk
			h2f_lw_AWID        => hps_0_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR      => hps_0_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN       => hps_0_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE      => hps_0_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST     => hps_0_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK      => hps_0_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE     => hps_0_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT      => hps_0_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID     => hps_0_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY     => hps_0_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID         => hps_0_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA       => hps_0_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB       => hps_0_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST       => hps_0_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID      => hps_0_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY      => hps_0_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID         => hps_0_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP       => hps_0_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID      => hps_0_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY      => hps_0_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID        => hps_0_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR      => hps_0_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN       => hps_0_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE      => hps_0_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST     => hps_0_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK      => hps_0_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE     => hps_0_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT      => hps_0_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID     => hps_0_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY     => hps_0_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID         => hps_0_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA       => hps_0_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP       => hps_0_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST       => hps_0_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID      => hps_0_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY      => hps_0_h2f_lw_axi_master_rready,  --                  .rready
			f2h_irq_p0         => hps_0_f2h_irq0_irq,              --          f2h_irq0.irq
			f2h_irq_p1         => hps_0_f2h_irq1_irq               --          f2h_irq1.irq
		);

	interrupt : component hps_interrupt
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_1_interrupt_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_interrupt_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_interrupt_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_interrupt_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_interrupt_s1_readdata,        --                    .readdata
			in_port    => open,                                           -- external_connection.export
			out_port   => open,                                           --                    .export
			irq        => irq_mapper_receiver0_irq                        --                 irq.irq
		);

	start : component hps_start
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_1_start_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_start_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_start_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_start_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_start_s1_readdata,        --                    .readdata
			in_port    => open,                                       -- external_connection.export
			out_port   => open                                        --                    .export
		);

	mm_interconnect_0 : component hps_mm_interconnect_0
		port map (
			hps_0_h2f_axi_master_awid                                        => hps_0_h2f_axi_master_awid,          --                                       hps_0_h2f_axi_master.awid
			hps_0_h2f_axi_master_awaddr                                      => hps_0_h2f_axi_master_awaddr,        --                                                           .awaddr
			hps_0_h2f_axi_master_awlen                                       => hps_0_h2f_axi_master_awlen,         --                                                           .awlen
			hps_0_h2f_axi_master_awsize                                      => hps_0_h2f_axi_master_awsize,        --                                                           .awsize
			hps_0_h2f_axi_master_awburst                                     => hps_0_h2f_axi_master_awburst,       --                                                           .awburst
			hps_0_h2f_axi_master_awlock                                      => hps_0_h2f_axi_master_awlock,        --                                                           .awlock
			hps_0_h2f_axi_master_awcache                                     => hps_0_h2f_axi_master_awcache,       --                                                           .awcache
			hps_0_h2f_axi_master_awprot                                      => hps_0_h2f_axi_master_awprot,        --                                                           .awprot
			hps_0_h2f_axi_master_awvalid                                     => hps_0_h2f_axi_master_awvalid,       --                                                           .awvalid
			hps_0_h2f_axi_master_awready                                     => hps_0_h2f_axi_master_awready,       --                                                           .awready
			hps_0_h2f_axi_master_wid                                         => hps_0_h2f_axi_master_wid,           --                                                           .wid
			hps_0_h2f_axi_master_wdata                                       => hps_0_h2f_axi_master_wdata,         --                                                           .wdata
			hps_0_h2f_axi_master_wstrb                                       => hps_0_h2f_axi_master_wstrb,         --                                                           .wstrb
			hps_0_h2f_axi_master_wlast                                       => hps_0_h2f_axi_master_wlast,         --                                                           .wlast
			hps_0_h2f_axi_master_wvalid                                      => hps_0_h2f_axi_master_wvalid,        --                                                           .wvalid
			hps_0_h2f_axi_master_wready                                      => hps_0_h2f_axi_master_wready,        --                                                           .wready
			hps_0_h2f_axi_master_bid                                         => hps_0_h2f_axi_master_bid,           --                                                           .bid
			hps_0_h2f_axi_master_bresp                                       => hps_0_h2f_axi_master_bresp,         --                                                           .bresp
			hps_0_h2f_axi_master_bvalid                                      => hps_0_h2f_axi_master_bvalid,        --                                                           .bvalid
			hps_0_h2f_axi_master_bready                                      => hps_0_h2f_axi_master_bready,        --                                                           .bready
			hps_0_h2f_axi_master_arid                                        => hps_0_h2f_axi_master_arid,          --                                                           .arid
			hps_0_h2f_axi_master_araddr                                      => hps_0_h2f_axi_master_araddr,        --                                                           .araddr
			hps_0_h2f_axi_master_arlen                                       => hps_0_h2f_axi_master_arlen,         --                                                           .arlen
			hps_0_h2f_axi_master_arsize                                      => hps_0_h2f_axi_master_arsize,        --                                                           .arsize
			hps_0_h2f_axi_master_arburst                                     => hps_0_h2f_axi_master_arburst,       --                                                           .arburst
			hps_0_h2f_axi_master_arlock                                      => hps_0_h2f_axi_master_arlock,        --                                                           .arlock
			hps_0_h2f_axi_master_arcache                                     => hps_0_h2f_axi_master_arcache,       --                                                           .arcache
			hps_0_h2f_axi_master_arprot                                      => hps_0_h2f_axi_master_arprot,        --                                                           .arprot
			hps_0_h2f_axi_master_arvalid                                     => hps_0_h2f_axi_master_arvalid,       --                                                           .arvalid
			hps_0_h2f_axi_master_arready                                     => hps_0_h2f_axi_master_arready,       --                                                           .arready
			hps_0_h2f_axi_master_rid                                         => hps_0_h2f_axi_master_rid,           --                                                           .rid
			hps_0_h2f_axi_master_rdata                                       => hps_0_h2f_axi_master_rdata,         --                                                           .rdata
			hps_0_h2f_axi_master_rresp                                       => hps_0_h2f_axi_master_rresp,         --                                                           .rresp
			hps_0_h2f_axi_master_rlast                                       => hps_0_h2f_axi_master_rlast,         --                                                           .rlast
			hps_0_h2f_axi_master_rvalid                                      => hps_0_h2f_axi_master_rvalid,        --                                                           .rvalid
			hps_0_h2f_axi_master_rready                                      => hps_0_h2f_axi_master_rready,        --                                                           .rready
			clk_0_clk_clk                                                    => clk_clk,                            --                                                  clk_0_clk.clk
			hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset, -- hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			K_reset1_reset_bridge_in_reset_reset                             => rst_controller_reset_out_reset,     --                             K_reset1_reset_bridge_in_reset.reset
			K_s1_address                                                     => mm_interconnect_0_k_s1_address,     --                                                       K_s1.address
			K_s1_write                                                       => mm_interconnect_0_k_s1_write,       --                                                           .write
			K_s1_readdata                                                    => mm_interconnect_0_k_s1_readdata,    --                                                           .readdata
			K_s1_writedata                                                   => mm_interconnect_0_k_s1_writedata,   --                                                           .writedata
			K_s1_byteenable                                                  => mm_interconnect_0_k_s1_byteenable,  --                                                           .byteenable
			K_s1_chipselect                                                  => mm_interconnect_0_k_s1_chipselect,  --                                                           .chipselect
			K_s1_clken                                                       => mm_interconnect_0_k_s1_clken,       --                                                           .clken
			M_s1_address                                                     => mm_interconnect_0_m_s1_address,     --                                                       M_s1.address
			M_s1_write                                                       => mm_interconnect_0_m_s1_write,       --                                                           .write
			M_s1_readdata                                                    => mm_interconnect_0_m_s1_readdata,    --                                                           .readdata
			M_s1_writedata                                                   => mm_interconnect_0_m_s1_writedata,   --                                                           .writedata
			M_s1_byteenable                                                  => mm_interconnect_0_m_s1_byteenable,  --                                                           .byteenable
			M_s1_chipselect                                                  => mm_interconnect_0_m_s1_chipselect,  --                                                           .chipselect
			M_s1_clken                                                       => mm_interconnect_0_m_s1_clken        --                                                           .clken
		);

	mm_interconnect_1 : component hps_mm_interconnect_1
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,              --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,            --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,             --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,            --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,           --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,            --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,           --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,            --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,           --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,           --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,               --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,             --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,             --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,             --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,            --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,            --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,               --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,             --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,            --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,            --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,              --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,            --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,             --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,            --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,           --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,            --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,           --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,            --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,           --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,           --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,               --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,             --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,             --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,             --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,            --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,            --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                   --                                                     clk_0_clk.clk
			CNT_N_reset_reset_bridge_in_reset_reset                             => rst_controller_reset_out_reset,            --                             CNT_N_reset_reset_bridge_in_reset.reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,        -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			a_s1_address                                                        => mm_interconnect_1_a_s1_address,            --                                                          a_s1.address
			a_s1_write                                                          => mm_interconnect_1_a_s1_write,              --                                                              .write
			a_s1_readdata                                                       => mm_interconnect_1_a_s1_readdata,           --                                                              .readdata
			a_s1_writedata                                                      => mm_interconnect_1_a_s1_writedata,          --                                                              .writedata
			a_s1_chipselect                                                     => mm_interconnect_1_a_s1_chipselect,         --                                                              .chipselect
			a_init_s1_address                                                   => mm_interconnect_1_a_init_s1_address,       --                                                     a_init_s1.address
			a_init_s1_write                                                     => mm_interconnect_1_a_init_s1_write,         --                                                              .write
			a_init_s1_readdata                                                  => mm_interconnect_1_a_init_s1_readdata,      --                                                              .readdata
			a_init_s1_writedata                                                 => mm_interconnect_1_a_init_s1_writedata,     --                                                              .writedata
			a_init_s1_chipselect                                                => mm_interconnect_1_a_init_s1_chipselect,    --                                                              .chipselect
			b_s1_address                                                        => mm_interconnect_1_b_s1_address,            --                                                          b_s1.address
			b_s1_write                                                          => mm_interconnect_1_b_s1_write,              --                                                              .write
			b_s1_readdata                                                       => mm_interconnect_1_b_s1_readdata,           --                                                              .readdata
			b_s1_writedata                                                      => mm_interconnect_1_b_s1_writedata,          --                                                              .writedata
			b_s1_chipselect                                                     => mm_interconnect_1_b_s1_chipselect,         --                                                              .chipselect
			b_init_s1_address                                                   => mm_interconnect_1_b_init_s1_address,       --                                                     b_init_s1.address
			b_init_s1_write                                                     => mm_interconnect_1_b_init_s1_write,         --                                                              .write
			b_init_s1_readdata                                                  => mm_interconnect_1_b_init_s1_readdata,      --                                                              .readdata
			b_init_s1_writedata                                                 => mm_interconnect_1_b_init_s1_writedata,     --                                                              .writedata
			b_init_s1_chipselect                                                => mm_interconnect_1_b_init_s1_chipselect,    --                                                              .chipselect
			c_s1_address                                                        => mm_interconnect_1_c_s1_address,            --                                                          c_s1.address
			c_s1_write                                                          => mm_interconnect_1_c_s1_write,              --                                                              .write
			c_s1_readdata                                                       => mm_interconnect_1_c_s1_readdata,           --                                                              .readdata
			c_s1_writedata                                                      => mm_interconnect_1_c_s1_writedata,          --                                                              .writedata
			c_s1_chipselect                                                     => mm_interconnect_1_c_s1_chipselect,         --                                                              .chipselect
			c_init_s1_address                                                   => mm_interconnect_1_c_init_s1_address,       --                                                     c_init_s1.address
			c_init_s1_write                                                     => mm_interconnect_1_c_init_s1_write,         --                                                              .write
			c_init_s1_readdata                                                  => mm_interconnect_1_c_init_s1_readdata,      --                                                              .readdata
			c_init_s1_writedata                                                 => mm_interconnect_1_c_init_s1_writedata,     --                                                              .writedata
			c_init_s1_chipselect                                                => mm_interconnect_1_c_init_s1_chipselect,    --                                                              .chipselect
			CNT_N_s1_address                                                    => mm_interconnect_1_cnt_n_s1_address,        --                                                      CNT_N_s1.address
			CNT_N_s1_write                                                      => mm_interconnect_1_cnt_n_s1_write,          --                                                              .write
			CNT_N_s1_readdata                                                   => mm_interconnect_1_cnt_n_s1_readdata,       --                                                              .readdata
			CNT_N_s1_writedata                                                  => mm_interconnect_1_cnt_n_s1_writedata,      --                                                              .writedata
			CNT_N_s1_chipselect                                                 => mm_interconnect_1_cnt_n_s1_chipselect,     --                                                              .chipselect
			d_s1_address                                                        => mm_interconnect_1_d_s1_address,            --                                                          d_s1.address
			d_s1_write                                                          => mm_interconnect_1_d_s1_write,              --                                                              .write
			d_s1_readdata                                                       => mm_interconnect_1_d_s1_readdata,           --                                                              .readdata
			d_s1_writedata                                                      => mm_interconnect_1_d_s1_writedata,          --                                                              .writedata
			d_s1_chipselect                                                     => mm_interconnect_1_d_s1_chipselect,         --                                                              .chipselect
			d_init_s1_address                                                   => mm_interconnect_1_d_init_s1_address,       --                                                     d_init_s1.address
			d_init_s1_write                                                     => mm_interconnect_1_d_init_s1_write,         --                                                              .write
			d_init_s1_readdata                                                  => mm_interconnect_1_d_init_s1_readdata,      --                                                              .readdata
			d_init_s1_writedata                                                 => mm_interconnect_1_d_init_s1_writedata,     --                                                              .writedata
			d_init_s1_chipselect                                                => mm_interconnect_1_d_init_s1_chipselect,    --                                                              .chipselect
			e_s1_address                                                        => mm_interconnect_1_e_s1_address,            --                                                          e_s1.address
			e_s1_write                                                          => mm_interconnect_1_e_s1_write,              --                                                              .write
			e_s1_readdata                                                       => mm_interconnect_1_e_s1_readdata,           --                                                              .readdata
			e_s1_writedata                                                      => mm_interconnect_1_e_s1_writedata,          --                                                              .writedata
			e_s1_chipselect                                                     => mm_interconnect_1_e_s1_chipselect,         --                                                              .chipselect
			e_init_s1_address                                                   => mm_interconnect_1_e_init_s1_address,       --                                                     e_init_s1.address
			e_init_s1_write                                                     => mm_interconnect_1_e_init_s1_write,         --                                                              .write
			e_init_s1_readdata                                                  => mm_interconnect_1_e_init_s1_readdata,      --                                                              .readdata
			e_init_s1_writedata                                                 => mm_interconnect_1_e_init_s1_writedata,     --                                                              .writedata
			e_init_s1_chipselect                                                => mm_interconnect_1_e_init_s1_chipselect,    --                                                              .chipselect
			f_s1_address                                                        => mm_interconnect_1_f_s1_address,            --                                                          f_s1.address
			f_s1_write                                                          => mm_interconnect_1_f_s1_write,              --                                                              .write
			f_s1_readdata                                                       => mm_interconnect_1_f_s1_readdata,           --                                                              .readdata
			f_s1_writedata                                                      => mm_interconnect_1_f_s1_writedata,          --                                                              .writedata
			f_s1_chipselect                                                     => mm_interconnect_1_f_s1_chipselect,         --                                                              .chipselect
			f_init_s1_address                                                   => mm_interconnect_1_f_init_s1_address,       --                                                     f_init_s1.address
			f_init_s1_write                                                     => mm_interconnect_1_f_init_s1_write,         --                                                              .write
			f_init_s1_readdata                                                  => mm_interconnect_1_f_init_s1_readdata,      --                                                              .readdata
			f_init_s1_writedata                                                 => mm_interconnect_1_f_init_s1_writedata,     --                                                              .writedata
			f_init_s1_chipselect                                                => mm_interconnect_1_f_init_s1_chipselect,    --                                                              .chipselect
			g_s1_address                                                        => mm_interconnect_1_g_s1_address,            --                                                          g_s1.address
			g_s1_write                                                          => mm_interconnect_1_g_s1_write,              --                                                              .write
			g_s1_readdata                                                       => mm_interconnect_1_g_s1_readdata,           --                                                              .readdata
			g_s1_writedata                                                      => mm_interconnect_1_g_s1_writedata,          --                                                              .writedata
			g_s1_chipselect                                                     => mm_interconnect_1_g_s1_chipselect,         --                                                              .chipselect
			g_init_s1_address                                                   => mm_interconnect_1_g_init_s1_address,       --                                                     g_init_s1.address
			g_init_s1_write                                                     => mm_interconnect_1_g_init_s1_write,         --                                                              .write
			g_init_s1_readdata                                                  => mm_interconnect_1_g_init_s1_readdata,      --                                                              .readdata
			g_init_s1_writedata                                                 => mm_interconnect_1_g_init_s1_writedata,     --                                                              .writedata
			g_init_s1_chipselect                                                => mm_interconnect_1_g_init_s1_chipselect,    --                                                              .chipselect
			h_s1_address                                                        => mm_interconnect_1_h_s1_address,            --                                                          h_s1.address
			h_s1_write                                                          => mm_interconnect_1_h_s1_write,              --                                                              .write
			h_s1_readdata                                                       => mm_interconnect_1_h_s1_readdata,           --                                                              .readdata
			h_s1_writedata                                                      => mm_interconnect_1_h_s1_writedata,          --                                                              .writedata
			h_s1_chipselect                                                     => mm_interconnect_1_h_s1_chipselect,         --                                                              .chipselect
			h_init_s1_address                                                   => mm_interconnect_1_h_init_s1_address,       --                                                     h_init_s1.address
			h_init_s1_write                                                     => mm_interconnect_1_h_init_s1_write,         --                                                              .write
			h_init_s1_readdata                                                  => mm_interconnect_1_h_init_s1_readdata,      --                                                              .readdata
			h_init_s1_writedata                                                 => mm_interconnect_1_h_init_s1_writedata,     --                                                              .writedata
			h_init_s1_chipselect                                                => mm_interconnect_1_h_init_s1_chipselect,    --                                                              .chipselect
			interrupt_s1_address                                                => mm_interconnect_1_interrupt_s1_address,    --                                                  interrupt_s1.address
			interrupt_s1_write                                                  => mm_interconnect_1_interrupt_s1_write,      --                                                              .write
			interrupt_s1_readdata                                               => mm_interconnect_1_interrupt_s1_readdata,   --                                                              .readdata
			interrupt_s1_writedata                                              => mm_interconnect_1_interrupt_s1_writedata,  --                                                              .writedata
			interrupt_s1_chipselect                                             => mm_interconnect_1_interrupt_s1_chipselect, --                                                              .chipselect
			start_s1_address                                                    => mm_interconnect_1_start_s1_address,        --                                                      start_s1.address
			start_s1_write                                                      => mm_interconnect_1_start_s1_write,          --                                                              .write
			start_s1_readdata                                                   => mm_interconnect_1_start_s1_readdata,       --                                                              .readdata
			start_s1_writedata                                                  => mm_interconnect_1_start_s1_writedata,      --                                                              .writedata
			start_s1_chipselect                                                 => mm_interconnect_1_start_s1_chipselect      --                                                              .chipselect
		);

	irq_mapper : component hps_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			sender_irq    => hps_0_f2h_irq0_irq        --    sender.irq
		);

	irq_mapper_001 : component hps_irq_mapper_001
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq1_irq  --    sender.irq
		);

	rst_controller : component hps_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component hps_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_1_cnt_n_s1_write_ports_inv <= not mm_interconnect_1_cnt_n_s1_write;

	mm_interconnect_1_a_init_s1_write_ports_inv <= not mm_interconnect_1_a_init_s1_write;

	mm_interconnect_1_b_init_s1_write_ports_inv <= not mm_interconnect_1_b_init_s1_write;

	mm_interconnect_1_c_init_s1_write_ports_inv <= not mm_interconnect_1_c_init_s1_write;

	mm_interconnect_1_d_init_s1_write_ports_inv <= not mm_interconnect_1_d_init_s1_write;

	mm_interconnect_1_e_init_s1_write_ports_inv <= not mm_interconnect_1_e_init_s1_write;

	mm_interconnect_1_f_init_s1_write_ports_inv <= not mm_interconnect_1_f_init_s1_write;

	mm_interconnect_1_g_init_s1_write_ports_inv <= not mm_interconnect_1_g_init_s1_write;

	mm_interconnect_1_h_init_s1_write_ports_inv <= not mm_interconnect_1_h_init_s1_write;

	mm_interconnect_1_a_s1_write_ports_inv <= not mm_interconnect_1_a_s1_write;

	mm_interconnect_1_b_s1_write_ports_inv <= not mm_interconnect_1_b_s1_write;

	mm_interconnect_1_c_s1_write_ports_inv <= not mm_interconnect_1_c_s1_write;

	mm_interconnect_1_d_s1_write_ports_inv <= not mm_interconnect_1_d_s1_write;

	mm_interconnect_1_e_s1_write_ports_inv <= not mm_interconnect_1_e_s1_write;

	mm_interconnect_1_f_s1_write_ports_inv <= not mm_interconnect_1_f_s1_write;

	mm_interconnect_1_g_s1_write_ports_inv <= not mm_interconnect_1_g_s1_write;

	mm_interconnect_1_h_s1_write_ports_inv <= not mm_interconnect_1_h_s1_write;

	mm_interconnect_1_start_s1_write_ports_inv <= not mm_interconnect_1_start_s1_write;

	mm_interconnect_1_interrupt_s1_write_ports_inv <= not mm_interconnect_1_interrupt_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of hps
